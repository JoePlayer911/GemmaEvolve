module TopModule (
    input [31:0] in,
    output [31:0] out
);

  // Write your code here
  assign out = 32'b0; // Place holder

endmodule
